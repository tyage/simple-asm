module P2;
endmodule