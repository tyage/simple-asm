module P1TEST;

endmodule